/////////////////////////////////////////////////////////////////////////
//                                                                     //
//   Modulename :  sys_defs.vh                                         //
//                                                                     //
//  Description :  This file has the macro-defines for macros used in  //
//                 the pipeline design.                                //
//                                                                     //
/////////////////////////////////////////////////////////////////////////


`ifndef __SYS_DEFS_VH__
`define __SYS_DEFS_VH__

//////////////////////////////////////////////
//
// final project definitions
//
// Revision 1 by Hanbo
// Added ARF, ROB, PRF, RS size definition 
//
// Revision 2 by Hanbo
// RF_FU_PACKET definition 

//
//////////////////////////////////////////////

`define ARF_SIZE 32					
`define ROB_SIZE 64						
`define PRF_SIZE 96
`define ARF_WIDTH $clog2(`ARF_SIZE)
`define ROB_WIDTH $clog2(`ROB_SIZE)
`define PRF_WIDTH $clog2(`PRF_SIZE)
`define RS_WIDTH $clog2(`RS_SIZE)
`define N_WAY 3
`define N_WIDTH 2
`define BTB_SIZE 16
`define BTB_WIDTH $clog2(`BTB_SIZE)
`define PHT_SIZE 8
`define PHT_WIDTH $clog2(`PHT_SIZE)
`define BHT_SIZE 8
`define BHT_WIDTH $clog2(`BHT_SIZE)
`define PREFET_SIZE 8
`define PREFET_WIDTH $clog2(`PREFET_SIZE)


//op_type+ready*2+prn*3+rob+imm+fu_type+pc+npc+use_prn*2+op1_select+op2_select+extra+inst
`define RS1_DATABUS_IN_WIDTH 5+2+(`PRF_WIDTH)*3+(`ROB_WIDTH)+(`IMM_WIDTH)+4+(`XLEN)+(`XLEN)+2+2+4+6+(`XLEN)
`define RS1_DATABUS_OUT_WIDTH 5+(`PRF_WIDTH)*3+(`ROB_WIDTH)+(`IMM_WIDTH)+4+(`XLEN)+(`XLEN)+2+2+4+4+(`XLEN)
`define RS_SIZE 16
`define IMM_WIDTH 32
`define FU_CNT 6
`define DATABUS_FU_ALLOC (`XLEN)*2+5+(`XLEN)*2+6+(`PRF_WIDTH)+(`IMM_WIDTH)+(`ROB_WIDTH)+(`XLEN)
`define CDB_DATABUS_OUT_WIDTH 3*(`XLEN)+(`PRF_WIDTH)+(`ROB_WIDTH)+4
`define DC_SIZE 32

`ifdef  SYNTH_TEST
`define DUT(mod) mod``_svsim
`else
`define DUT(mod) mod
`endif

//////////////////////////////////////////////
//
// Memory/testbench attribute definitions
//
//////////////////////////////////////////////
`define CACHE_MODE //removes the byte-level interface from the memory mode, DO NOT MODIFY!
`define NUM_MEM_TAGS           15 //num of outstanding requests the memory can handle

`define MEM_SIZE_IN_BYTES      (64*1024)
`define MEM_64BIT_LINES        (`MEM_SIZE_IN_BYTES/8)

//you can change the clock period to whatever, 10 is just fine
`define VERILOG_CLOCK_PERIOD   10.0
`define SYNTH_CLOCK_PERIOD     10.0 // Clock period for synth and memory latency

`define MEM_LATENCY_IN_CYCLES (100.0/`SYNTH_CLOCK_PERIOD+0.49999)
// the 0.49999 is to force ceiling(100/period).  The default behavior for
// float to integer conversion is rounding to nearest

typedef union packed {
    logic [7:0][7:0] byte_level;
    logic [3:0][15:0] half_level;
    logic [1:0][31:0] word_level;
} EXAMPLE_CACHE_BLOCK;

//////////////////////////////////////////////
// Exception codes
// This mostly follows the RISC-V Privileged spec
// except a few add-ons for our infrastructure
// The majority of them won't be used, but it's
// good to know what they are
//////////////////////////////////////////////

typedef enum logic [3:0] {
	INST_ADDR_MISALIGN  = 4'h0,
	INST_ACCESS_FAULT   = 4'h1,
	ILLEGAL_INST        = 4'h2,
	BREAKPOINT          = 4'h3,
	LOAD_ADDR_MISALIGN  = 4'h4,
	LOAD_ACCESS_FAULT   = 4'h5,
	STORE_ADDR_MISALIGN = 4'h6,
	STORE_ACCESS_FAULT  = 4'h7,
	ECALL_U_MODE        = 4'h8,
	ECALL_S_MODE        = 4'h9,
	NO_ERROR            = 4'ha, //a reserved code that we modified for our purpose
	ECALL_M_MODE        = 4'hb,
	INST_PAGE_FAULT     = 4'hc,
	LOAD_PAGE_FAULT     = 4'hd,
	HALTED_ON_WFI       = 4'he, //another reserved code that we used
	STORE_PAGE_FAULT    = 4'hf
} EXCEPTION_CODE;


//////////////////////////////////////////////
//
// Datapath control signals
//
//////////////////////////////////////////////

//
// ALU opA input mux selects
//
typedef enum logic [1:0] {
	OPA_IS_RS1  = 2'h0,
	OPA_IS_NPC  = 2'h1,
	OPA_IS_PC   = 2'h2,
	OPA_IS_ZERO = 2'h3
} ALU_OPA_SELECT;

//
// ALU opB input mux selects
//
typedef enum logic [3:0] {
	OPB_IS_RS2    = 4'h0,
	OPB_IS_I_IMM  = 4'h1,
	OPB_IS_S_IMM  = 4'h2,
	OPB_IS_B_IMM  = 4'h3,
	OPB_IS_U_IMM  = 4'h4,
	OPB_IS_J_IMM  = 4'h5
} ALU_OPB_SELECT;

//
// Destination register select
//
typedef enum logic [1:0] {
	DEST_RD = 2'h0,
	DEST_NONE  = 2'h1
} DEST_REG_SEL;

//
// ALU function code input
// probably want to leave these alone
//
typedef enum logic [4:0] {
	ALU_ADD     = 5'h00,
	ALU_SUB     = 5'h01,
	ALU_SLT     = 5'h02,
	ALU_SLTU    = 5'h03,
	ALU_AND     = 5'h04,
	ALU_OR      = 5'h05,
	ALU_XOR     = 5'h06,
	ALU_SLL     = 5'h07,
	ALU_SRL     = 5'h08,
	ALU_SRA     = 5'h09,
	ALU_MUL     = 5'h0a,
	ALU_MULH    = 5'h0b,
	ALU_MULHSU  = 5'h0c,
	ALU_MULHU   = 5'h0d,
	ALU_DIV     = 5'h0e,
	ALU_DIVU    = 5'h0f,
	ALU_REM     = 5'h10,
	ALU_REMU    = 5'h11
} ALU_FUNC;

//////////////////////////////////////////////
//
// Assorted things it is not wise to change
//
//////////////////////////////////////////////

//
// actually, you might have to change this if you change VERILOG_CLOCK_PERIOD
// JK you don't ^^^
//
`define SD #1


// the RISCV register file zero register, any read of this register always
// returns a zero value, and any write to this register is thrown away
//
`define ZERO_REG 5'd0

//
// Memory bus commands control signals
//
typedef enum logic [1:0] {
	BUS_NONE     = 2'h0,
	BUS_LOAD     = 2'h1,
	BUS_STORE    = 2'h2
} BUS_COMMAND;


typedef enum logic [1:0] {
	BYTE = 2'h0,
	HALF = 2'h1,
	WORD = 2'h2,
	DOUBLE = 2'h3
} MEM_SIZE;

//
// useful boolean single-bit definitions
//
`define FALSE  1'h0
`define TRUE  1'h1

// RISCV ISA SPEC
`define XLEN 32
typedef union packed {
	logic [31:0] inst;
	struct packed {
		logic [6:0] funct7;
		logic [4:0] rs2;
		logic [4:0] rs1;
		logic [2:0] funct3;
		logic [4:0] rd;
		logic [6:0] opcode;
	} r; //register to register instructions
	struct packed {
		logic [11:0] imm;
		logic [4:0]  rs1; //base
		logic [2:0]  funct3;
		logic [4:0]  rd;  //dest
		logic [6:0]  opcode;
	} i; //immediate or load instructions
	struct packed {
		logic [6:0] off; //offset[11:5] for calculating address
		logic [4:0] rs2; //source
		logic [4:0] rs1; //base
		logic [2:0] funct3;
		logic [4:0] set; //offset[4:0] for calculating address
		logic [6:0] opcode;
	} s; //store instructions
	struct packed {
		logic       of; //offset[12]
		logic [5:0] s;   //offset[10:5]
		logic [4:0] rs2;//source 2
		logic [4:0] rs1;//source 1
		logic [2:0] funct3;
		logic [3:0] et; //offset[4:1]
		logic       f;  //offset[11]
		logic [6:0] opcode;
	} b; //branch instructions
	struct packed {
		logic [19:0] imm;
		logic [4:0]  rd;
		logic [6:0]  opcode;
	} u; //upper immediate instructions
	struct packed {
		logic       of; //offset[20]
		logic [9:0] et; //offset[10:1]
		logic       s;  //offset[11]
		logic [7:0] f;	//offset[19:12]
		logic [4:0] rd; //dest
		logic [6:0] opcode;
	} j;  //jump instructions
`ifdef ATOMIC_EXT
	struct packed {
		logic [4:0] funct5;
		logic       aq;
		logic       rl;
		logic [4:0] rs2;
		logic [4:0] rs1;
		logic [2:0] funct3;
		logic [4:0] rd;
		logic [6:0] opcode;
	} a; //atomic instructions
`endif
`ifdef SYSTEM_EXT
	struct packed {
		logic [11:0] csr;
		logic [4:0]  rs1;
		logic [2:0]  funct3;
		logic [4:0]  rd;
		logic [6:0]  opcode;
	} sys; //system call instructions
`endif

} INST; //instruction typedef, this should cover all types of instructions

//
// Basic NOP instruction.  Allows pipline registers to clearly be reset with
// an instruction that does nothing instead of Zero which is really an ADDI x0, x0, 0
//
`define NOP 32'h00000013

//////////////////////////////////////////////
//
// IF Packets:
// Data that is exchanged between the IF and the ID stages  
//
//////////////////////////////////////////////
typedef struct packed {
	logic uncond_branch;			// if the branch is unconditional
        logic cond_branch;			// if the branch is conditional
////////Predictor outputs
	logic branch_is_taken;			// is branch predicted taken/not taken? (by local predictor)
	logic [`XLEN-1:0] branch_PC;		// the PC for the branch
	logic [`XLEN-1:0] branch_target_PC;	// the target address by BTB
////////FU outputs
	logic branch_true_taken;		// is the brach actually taken? (calculated by FU)
	logic [`XLEN-1:0] branch_true_target_PC;// the true target address for the branch (calculated by FU)
////////Misprediction (ROB commit outputs)
	logic branch_misprediction;		// If the branch is mispredicted
	logic [`XLEN-1:0] branch_true_PC;	// The true target PC after misprediction	
} ROB_IF_BRANCH_PACKET;

typedef struct packed {
	logic valid; 					// If low, the data in this struct is garbage
        INST  inst; 					// fetched instruction out
	logic [`XLEN-1:0] NPC; 				// PC + 4
	logic [`XLEN-1:0] PC;  				// PC 
	logic	   	  branch_predicted_taken; 	// From predictor, indicating if the branch is taken/not taken
	logic [`XLEN-1:0] branch_predicted_PC;    	// The predicted target PC from predictor	
} IF_ID_PACKET;

//////////////////////////////////////////////
//
// ID Packets:
// Data that is exchanged from ID to EX stage
//
//////////////////////////////////////////////

typedef struct packed {
	logic [`XLEN-1:0] NPC;   // PC + 4
	logic [`XLEN-1:0] PC;    // PC

	logic [3:0]	  FU_type; 		 // branch,mem,mul,alu
	logic [`PRF_WIDTH-1:0] rs1_prf_value;    // reg A prf value  
	logic		  rs1_use_prf;		 // if reg A prf is needed
	logic		  rs1_prf_valid;	 // is rs1_prf valid                               
	logic [`XLEN-1:0] rs1_nprf_value;	 // Operand A is PC or NPC
	logic		  rs1_is_nprf;		 // is opa not prf
	logic [`PRF_WIDTH-1:0] rs2_prf_value;    // reg B prf value  
	logic		  rs2_use_prf;		 // if reg B prf is needed 
	logic		  rs2_prf_valid;      	 // is rs2_prf valid         
	logic [`XLEN-1:0] rs2_nprf_value;	 // Operand B is immediate
	logic		  rs2_is_imm;    	 // is opb an immediate              
	                                                                                
	ALU_OPA_SELECT opa_select; 		// ALU opa mux select (ALU_OPA_xxx *)
	ALU_OPB_SELECT opb_select; 		// ALU opb mux select (ALU_OPB_xxx *)
	INST inst;                 		// instruction
	
	logic [4:0] dest_reg_idx;  		// destination (writeback) register arf index    
	logic [`PRF_WIDTH-1:0] dest_prf_reg; 	// destination register prf index
	logic [`PRF_WIDTH-1:0] dest_old_prn; 	// old prn value of the destination register
	ALU_FUNC    alu_func;      		// ALU function select (ALU_xxx *)
	logic       rd_mem;        		// does inst read memory?
	logic       wr_mem;        		// does inst write memory?
	logic       cond_branch;   		// is inst a conditional branch?
	logic       uncond_branch; 		// is inst an unconditional branch?
	logic	    branch_predict;		//taken/not taken
	logic [`XLEN-1:0]	predict_PC;
	logic       halt;          		// is this a halt?
	logic       illegal;       		// is this instruction illegal?
	logic       csr_op;       		// is this a CSR operation? (we only used this as a cheap way to get return code)
	logic       valid;        		// is inst a valid instruction to be counted for CPI calculations?
} ID_EX_PACKET;

typedef struct packed {
	logic [`XLEN-1:0] alu_result; 		// alu_result
	logic [`XLEN-1:0] NPC; 			//pc + 4
	logic             take_branch; 		// is this a taken branch?
	//pass throughs from decode stage
	logic [`XLEN-1:0] rs2_value;
	logic             rd_mem, wr_mem;
	logic [4:0]       dest_reg_idx;
	logic             halt, illegal, csr_op, valid;
	logic [2:0]       mem_size; 		// byte, half-word or word
} EX_MEM_PACKET;

typedef struct packed {
	logic		  	valid;
	logic		  	commit; 		// 0: not yet executed,1 execution finish(by CDB)
	logic 			branch_true_taken;	// is the brach actually taken? (calculated by FU)
	logic [`XLEN-1:0] 	branch_true_target_PC;	// the true target address for the branch (calculated by FU)
	logic		  	branch_mispredict;
	logic [`XLEN-1:0] 	branch_true_PC;		// The true PC after misprediction
	logic [`XLEN-1:0] 	proc2mem_addr;     	// Address sent to memory
	logic [63:0] 		proc2mem_data;      	// Data sent to memory
	logic [2:0] 		proc2mem_size;          // data size sent to memory
	ID_EX_PACKET 		id_packet;
} ROB_PACKET;

typedef struct packed {
	logic		  	valid;			//if this is a valid request
	logic		  	send; 			//if this request is sent to memory
	logic [3:0]		mem_tag;		//the tag derived from memory
	logic [`XLEN-1:0]	addr;			//the address of the request
	logic [4:0]		idx;			//the index of the request address
	logic [7:0] 		tag;			//the tag of the reqeust address
	logic [63:0] 		data;			//the data get from the memory
	logic			write_en;		//already get the data and ready to be writen to memory
} PREFETCHER_PACKET;


`endif // __SYS_DEFS_VH__
